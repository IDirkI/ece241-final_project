`timescale 1ns / 1ps

module testbench ( );

	parameter WOI = 9;
	parameter WOF = 16;

	wire [2:0][3:0][WOI+WOF-1:0] Poly1;
	wire [2:0][3:0][WOI+WOF-1:0] Poly2;
	wire [2:0][3:0][WOI+WOF-1:0] Poly3;
	wire [2:0][3:0][WOI+WOF-1:0] Poly4;
	wire [2:0][3:0][WOI+WOF-1:0] Poly5;
	wire [2:0][3:0][WOI+WOF-1:0] Poly6;
	wire [2:0][3:0][WOI+WOF-1:0] Poly7;
	wire [2:0][3:0][WOI+WOF-1:0] Poly8;
	wire [2:0][3:0][WOI+WOF-1:0] Poly9;
	wire [2:0][3:0][WOI+WOF-1:0] Poly10;
	wire [2:0][3:0][WOI+WOF-1:0] Poly11;
	wire [2:0][3:0][WOI+WOF-1:0] Poly12;
	
	initial begin
	end // initial
	Polygon_List U1 (Poly1, Poly2, Poly3, Poly4, Poly5, Poly6, Poly7, Poly8, Poly9, Poly10, Poly11, Poly12);

endmodule
