module Projector # (
		parameter	WII = 9,
						WIF = 16,
						WOI = 9,
						WOF = 16
		) (	
		// Inputs
			position,
			orientation,
			Polygon_in,
		// Outputs
			Polygon_out
);
/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/
 
/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
 // Inputs
 input wire 	signed 	[2:0][WOI+WOF-1:0] position;
 input wire 	signed 	[2:0][WOI+WOF-1:0] orientation;
 input wire 	signed 	[2:0][3:0][WII+WIF-1:0] Polygon_in;
 
 // Bidirectionals
 inout logic 	signed	[2:0][3:0][WII+WIF-1:0] Polygon_out;
	
/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
 
/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/

/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/
 
/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/
 projection # (
	.WII(WII), .WIF(WIF),
	.WOI(WOI), .WOF(WOF)
	) proj (.position(position), .orientation(orientation), .Polygon_in(Polygon_in), .Polygon_out(Polygon_out));
	

endmodule
